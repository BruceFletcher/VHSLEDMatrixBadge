library verilog;
use verilog.vl_types.all;
entity shhh_5th_cpld_tb is
end shhh_5th_cpld_tb;
